//------------------------------------------------------------------------------
// File       : opcodes.sv
// Author     : Lewis Russell
// Description: Definition of opcodes for picomips instructions set.
//------------------------------------------------------------------------------
parameter OP_LSW  = 6'b000110;
parameter OP_RTA  = 6'b000000;
parameter OP_ATR  = 6'b010111;
parameter OP_ADD  = 6'b000001;
parameter OP_ADDI = 6'b000101;
parameter OP_MULI = 6'b001011;
parameter OP_HEI  = 6'b100100;
