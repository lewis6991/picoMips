//------------------------------------------------------------------------------
// File       : opcodes.sv
// Author     : Lewis Russell
// Description: Definition of opcodes for picomips instructions set.
//------------------------------------------------------------------------------
parameter OP_LSW  = 7'b0000010;
parameter OP_RTA  = 7'b1000000;
parameter OP_ATR  = 7'b0010001;
parameter OP_ADD  = 7'b1000001;
parameter OP_ADDI = 7'b0000101;
parameter OP_MULI = 7'b0001011;
parameter OP_HEI  = 7'b0100100;
