//------------------------------------------------------------------------------
// File       : opcodes.sv
// Author     : Lewis Russell
// Description: Definition of opcodes for picomips instructions set.
//------------------------------------------------------------------------------
parameter OP_LSW  = 3'b110;
parameter OP_RTA  = 3'b000;
parameter OP_ATR  = 3'b111;
parameter OP_ADD  = 3'b001;
parameter OP_ADDI = 3'b101;
parameter OP_MULI = 3'b011;
parameter OP_HEI  = 3'b100;
