//------------------------------------------------------------------------------
// File       : opcodes.sv
// Author     : Lewis Russell
// Description: Definition of opcodes for picomips instructions set.
//------------------------------------------------------------------------------
parameter OP_LSW  = 6'b000010;
parameter OP_RTA  = 6'b100000;
parameter OP_ATR  = 6'b001001;
parameter OP_ADD  = 6'b100001;
parameter OP_ADDI = 6'b000101;
parameter OP_MULI = 6'b000001;
parameter OP_HEI  = 6'b010100;
